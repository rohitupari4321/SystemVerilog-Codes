interface intf();
  
  logic [3:0]i;
  logic [1:0]s;
  logic y;
  
  // interface also contains clocking block and mod port they aren't used here as it isn't a big design.
  
endinterface
interface intf();
  
  logic a;
  logic b;
  logic sum;
  logic carry;
  
  // interface also contains clocking block and mod port they aren't used here as it isn't a big design.
  
endinterface